module and_op (a, b, c);
  // a
  `include "included.svh"
endmodule
