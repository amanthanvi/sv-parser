/* IEEE1800-2017 Clause 22.5.1 page 680
*/

`define append(f) f``_master

module clock_master;
endmodule
