module A;
wire a = 1'b0;


endmodule
