module and_op (a, b, c);
 
endmodule
