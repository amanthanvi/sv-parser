module and_op (a, b, c);
`include "included.svh"   `include "included.svh"
endmodule
