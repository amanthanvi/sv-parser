`define PATH "included.svh"
module and_op (a, b, c);
`include `PATH
endmodule
