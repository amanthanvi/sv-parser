module and_op (a, b, c);
`include "included.svh" endmodule
