`define PATH included.svh
`define QUOTED_PATH `"`PATH`"
module and_op (a, b, c);
`include `QUOTED_PATH
endmodule
