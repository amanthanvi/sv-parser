`ifndef X
// pragma translate_off
module A;
endmodule
// pragma translate_on
`endif
