`define b `c
`define c `d
`define d `e
`define e `b
// indirect recursion
`b
