// foo
`include "include_recursive.svh"
// bar
